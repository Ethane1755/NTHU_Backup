module not_gate (
    input a,
    output o
);

not (o, a);

endmodule

module and_gate (
    input a,
    input b,
    output o1
);

and (o1, a, b);

endmodule


